** sch_path: /home/nvm_user4/RRAM_IMC/xschem/user_analog_project_wrapper.sch
.subckt user_analog_project_wrapper vdda1 vdda2 vssa1 vssa2 vccd1 vccd2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_stb_i wbs_cyc_i wbs_we_i wbs_sel_i[3] wbs_sel_i[2] wbs_sel_i[1] wbs_sel_i[0] wbs_dat_i[31]
+ wbs_dat_i[30] wbs_dat_i[29] wbs_dat_i[28] wbs_dat_i[27] wbs_dat_i[26] wbs_dat_i[25] wbs_dat_i[24] wbs_dat_i[23]
+ wbs_dat_i[22] wbs_dat_i[21] wbs_dat_i[20] wbs_dat_i[19] wbs_dat_i[18] wbs_dat_i[17] wbs_dat_i[16] wbs_dat_i[15]
+ wbs_dat_i[14] wbs_dat_i[13] wbs_dat_i[12] wbs_dat_i[11] wbs_dat_i[10] wbs_dat_i[9] wbs_dat_i[8] wbs_dat_i[7]
+ wbs_dat_i[6] wbs_dat_i[5] wbs_dat_i[4] wbs_dat_i[3] wbs_dat_i[2] wbs_dat_i[1] wbs_dat_i[0] wbs_adr_i[31]
+ wbs_adr_i[30] wbs_adr_i[29] wbs_adr_i[28] wbs_adr_i[27] wbs_adr_i[26] wbs_adr_i[25] wbs_adr_i[24] wbs_adr_i[23]
+ wbs_adr_i[22] wbs_adr_i[21] wbs_adr_i[20] wbs_adr_i[19] wbs_adr_i[18] wbs_adr_i[17] wbs_adr_i[16] wbs_adr_i[15]
+ wbs_adr_i[14] wbs_adr_i[13] wbs_adr_i[12] wbs_adr_i[11] wbs_adr_i[10] wbs_adr_i[9] wbs_adr_i[8] wbs_adr_i[7]
+ wbs_adr_i[6] wbs_adr_i[5] wbs_adr_i[4] wbs_adr_i[3] wbs_adr_i[2] wbs_adr_i[1] wbs_adr_i[0] wbs_ack_o
+ wbs_dat_o[31] wbs_dat_o[30] wbs_dat_o[29] wbs_dat_o[28] wbs_dat_o[27] wbs_dat_o[26] wbs_dat_o[25] wbs_dat_o[24]
+ wbs_dat_o[23] wbs_dat_o[22] wbs_dat_o[21] wbs_dat_o[20] wbs_dat_o[19] wbs_dat_o[18] wbs_dat_o[17] wbs_dat_o[16]
+ wbs_dat_o[15] wbs_dat_o[14] wbs_dat_o[13] wbs_dat_o[12] wbs_dat_o[11] wbs_dat_o[10] wbs_dat_o[9] wbs_dat_o[8]
+ wbs_dat_o[7] wbs_dat_o[6] wbs_dat_o[5] wbs_dat_o[4] wbs_dat_o[3] wbs_dat_o[2] wbs_dat_o[1] wbs_dat_o[0]
+ la_data_in[127] la_data_in[126] la_data_in[125] la_data_in[124] la_data_in[123] la_data_in[122] la_data_in[121]
+ la_data_in[120] la_data_in[119] la_data_in[118] la_data_in[117] la_data_in[116] la_data_in[115] la_data_in[114]
+ la_data_in[113] la_data_in[112] la_data_in[111] la_data_in[110] la_data_in[109] la_data_in[108] la_data_in[107]
+ la_data_in[106] la_data_in[105] la_data_in[104] la_data_in[103] la_data_in[102] la_data_in[101] la_data_in[100]
+ la_data_in[99] la_data_in[98] la_data_in[97] la_data_in[96] la_data_in[95] la_data_in[94] la_data_in[93]
+ la_data_in[92] la_data_in[91] la_data_in[90] la_data_in[89] la_data_in[88] la_data_in[87] la_data_in[86]
+ la_data_in[85] la_data_in[84] la_data_in[83] la_data_in[82] la_data_in[81] la_data_in[80] la_data_in[79]
+ la_data_in[78] la_data_in[77] la_data_in[76] la_data_in[75] la_data_in[74] la_data_in[73] la_data_in[72]
+ la_data_in[71] la_data_in[70] la_data_in[69] la_data_in[68] la_data_in[67] la_data_in[66] la_data_in[65]
+ la_data_in[64] la_data_in[63] la_data_in[62] la_data_in[61] la_data_in[60] la_data_in[59] la_data_in[58]
+ la_data_in[57] la_data_in[56] la_data_in[55] la_data_in[54] la_data_in[53] la_data_in[52] la_data_in[51]
+ la_data_in[50] la_data_in[49] la_data_in[48] la_data_in[47] la_data_in[46] la_data_in[45] la_data_in[44]
+ la_data_in[43] la_data_in[42] la_data_in[41] la_data_in[40] la_data_in[39] la_data_in[38] la_data_in[37]
+ la_data_in[36] la_data_in[35] la_data_in[34] la_data_in[33] la_data_in[32] la_data_in[31] la_data_in[30]
+ la_data_in[29] la_data_in[28] la_data_in[27] la_data_in[26] la_data_in[25] la_data_in[24] la_data_in[23]
+ la_data_in[22] la_data_in[21] la_data_in[20] la_data_in[19] la_data_in[18] la_data_in[17] la_data_in[16]
+ la_data_in[15] la_data_in[14] la_data_in[13] la_data_in[12] la_data_in[11] la_data_in[10] la_data_in[9]
+ la_data_in[8] la_data_in[7] la_data_in[6] la_data_in[5] la_data_in[4] la_data_in[3] la_data_in[2] la_data_in[1]
+ la_data_in[0] la_data_out[127] la_data_out[126] la_data_out[125] la_data_out[124] la_data_out[123]
+ la_data_out[122] la_data_out[121] la_data_out[120] la_data_out[119] la_data_out[118] la_data_out[117]
+ la_data_out[116] la_data_out[115] la_data_out[114] la_data_out[113] la_data_out[112] la_data_out[111]
+ la_data_out[110] la_data_out[109] la_data_out[108] la_data_out[107] la_data_out[106] la_data_out[105]
+ la_data_out[104] la_data_out[103] la_data_out[102] la_data_out[101] la_data_out[100] la_data_out[99] la_data_out[98]
+ la_data_out[97] la_data_out[96] la_data_out[95] la_data_out[94] la_data_out[93] la_data_out[92] la_data_out[91]
+ la_data_out[90] la_data_out[89] la_data_out[88] la_data_out[87] la_data_out[86] la_data_out[85] la_data_out[84]
+ la_data_out[83] la_data_out[82] la_data_out[81] la_data_out[80] la_data_out[79] la_data_out[78] la_data_out[77]
+ la_data_out[76] la_data_out[75] la_data_out[74] la_data_out[73] la_data_out[72] la_data_out[71] la_data_out[70]
+ la_data_out[69] la_data_out[68] la_data_out[67] la_data_out[66] la_data_out[65] la_data_out[64] la_data_out[63]
+ la_data_out[62] la_data_out[61] la_data_out[60] la_data_out[59] la_data_out[58] la_data_out[57] la_data_out[56]
+ la_data_out[55] la_data_out[54] la_data_out[53] la_data_out[52] la_data_out[51] la_data_out[50] la_data_out[49]
+ la_data_out[48] la_data_out[47] la_data_out[46] la_data_out[45] la_data_out[44] la_data_out[43] la_data_out[42]
+ la_data_out[41] la_data_out[40] la_data_out[39] la_data_out[38] la_data_out[37] la_data_out[36] la_data_out[35]
+ la_data_out[34] la_data_out[33] la_data_out[32] la_data_out[31] la_data_out[30] la_data_out[29] la_data_out[28]
+ la_data_out[27] la_data_out[26] la_data_out[25] la_data_out[24] la_data_out[23] la_data_out[22] la_data_out[21]
+ la_data_out[20] la_data_out[19] la_data_out[18] la_data_out[17] la_data_out[16] la_data_out[15] la_data_out[14]
+ la_data_out[13] la_data_out[12] la_data_out[11] la_data_out[10] la_data_out[9] la_data_out[8] la_data_out[7]
+ la_data_out[6] la_data_out[5] la_data_out[4] la_data_out[3] la_data_out[2] la_data_out[1] la_data_out[0] io_in[26]
+ io_in[25] io_in[24] io_in[23] io_in[22] io_in[21] io_in[20] io_in[19] io_in[18] io_in[17] io_in[16] io_in[15]
+ io_in[14] io_in[13] io_in[12] io_in[11] io_in[10] io_in[9] io_in[8] io_in[7] io_in[6] io_in[5] io_in[4]
+ io_in[3] io_in[2] io_in[1] io_in[0] io_in_3v3[26] io_in_3v3[25] io_in_3v3[24] io_in_3v3[23] io_in_3v3[22]
+ io_in_3v3[21] io_in_3v3[20] io_in_3v3[19] io_in_3v3[18] io_in_3v3[17] io_in_3v3[16] io_in_3v3[15] io_in_3v3[14]
+ io_in_3v3[13] io_in_3v3[12] io_in_3v3[11] io_in_3v3[10] io_in_3v3[9] io_in_3v3[8] io_in_3v3[7] io_in_3v3[6]
+ io_in_3v3[5] io_in_3v3[4] io_in_3v3[3] io_in_3v3[2] io_in_3v3[1] io_in_3v3[0] user_clock2 io_out[26] io_out[25]
+ io_out[24] io_out[23] io_out[22] io_out[21] io_out[20] io_out[19] io_out[18] io_out[17] io_out[16] io_out[15]
+ io_out[14] io_out[13] io_out[12] io_out[11] io_out[10] io_out[9] io_out[8] io_out[7] io_out[6] io_out[5]
+ io_out[4] io_out[3] io_out[2] io_out[1] io_out[0] io_oeb[26] io_oeb[25] io_oeb[24] io_oeb[23] io_oeb[22]
+ io_oeb[21] io_oeb[20] io_oeb[19] io_oeb[18] io_oeb[17] io_oeb[16] io_oeb[15] io_oeb[14] io_oeb[13] io_oeb[12]
+ io_oeb[11] io_oeb[10] io_oeb[9] io_oeb[8] io_oeb[7] io_oeb[6] io_oeb[5] io_oeb[4] io_oeb[3] io_oeb[2]
+ io_oeb[1] io_oeb[0] gpio_analog[17] gpio_analog[16] gpio_analog[15] gpio_analog[14] gpio_analog[13]
+ gpio_analog[12] gpio_analog[11] gpio_analog[10] gpio_analog[9] gpio_analog[8] gpio_analog[7] gpio_analog[6]
+ gpio_analog[5] gpio_analog[4] gpio_analog[3] gpio_analog[2] gpio_analog[1] gpio_analog[0] gpio_noesd[17]
+ gpio_noesd[16] gpio_noesd[15] gpio_noesd[14] gpio_noesd[13] gpio_noesd[12] gpio_noesd[11] gpio_noesd[10]
+ gpio_noesd[9] gpio_noesd[8] gpio_noesd[7] gpio_noesd[6] gpio_noesd[5] gpio_noesd[4] gpio_noesd[3] gpio_noesd[2]
+ gpio_noesd[1] gpio_noesd[0] io_analog[10] io_analog[9] io_analog[8] io_analog[7] io_analog[6] io_analog[5]
+ io_analog[4] io_analog[3] io_analog[2] io_analog[1] io_analog[0] io_clamp_high[2] io_clamp_high[1]
+ io_clamp_high[0] io_clamp_low[2] io_clamp_low[1] io_clamp_low[0] user_irq[2] user_irq[1] user_irq[0] la_oenb[127]
+ la_oenb[126] la_oenb[125] la_oenb[124] la_oenb[123] la_oenb[122] la_oenb[121] la_oenb[120] la_oenb[119]
+ la_oenb[118] la_oenb[117] la_oenb[116] la_oenb[115] la_oenb[114] la_oenb[113] la_oenb[112] la_oenb[111]
+ la_oenb[110] la_oenb[109] la_oenb[108] la_oenb[107] la_oenb[106] la_oenb[105] la_oenb[104] la_oenb[103]
+ la_oenb[102] la_oenb[101] la_oenb[100] la_oenb[99] la_oenb[98] la_oenb[97] la_oenb[96] la_oenb[95] la_oenb[94]
+ la_oenb[93] la_oenb[92] la_oenb[91] la_oenb[90] la_oenb[89] la_oenb[88] la_oenb[87] la_oenb[86] la_oenb[85]
+ la_oenb[84] la_oenb[83] la_oenb[82] la_oenb[81] la_oenb[80] la_oenb[79] la_oenb[78] la_oenb[77] la_oenb[76]
+ la_oenb[75] la_oenb[74] la_oenb[73] la_oenb[72] la_oenb[71] la_oenb[70] la_oenb[69] la_oenb[68] la_oenb[67]
+ la_oenb[66] la_oenb[65] la_oenb[64] la_oenb[63] la_oenb[62] la_oenb[61] la_oenb[60] la_oenb[59] la_oenb[58]
+ la_oenb[57] la_oenb[56] la_oenb[55] la_oenb[54] la_oenb[53] la_oenb[52] la_oenb[51] la_oenb[50] la_oenb[49]
+ la_oenb[48] la_oenb[47] la_oenb[46] la_oenb[45] la_oenb[44] la_oenb[43] la_oenb[42] la_oenb[41] la_oenb[40]
+ la_oenb[39] la_oenb[38] la_oenb[37] la_oenb[36] la_oenb[35] la_oenb[34] la_oenb[33] la_oenb[32] la_oenb[31]
+ la_oenb[30] la_oenb[29] la_oenb[28] la_oenb[27] la_oenb[26] la_oenb[25] la_oenb[24] la_oenb[23] la_oenb[22]
+ la_oenb[21] la_oenb[20] la_oenb[19] la_oenb[18] la_oenb[17] la_oenb[16] la_oenb[15] la_oenb[14] la_oenb[13]
+ la_oenb[12] la_oenb[11] la_oenb[10] la_oenb[9] la_oenb[8] la_oenb[7] la_oenb[6] la_oenb[5] la_oenb[4]
+ la_oenb[3] la_oenb[2] la_oenb[1] la_oenb[0]
*.PININFO vdda1:B vdda2:B vssa1:B vssa2:B vccd1:B vccd2:B vssd1:B vssd2:B wb_clk_i:I wb_rst_i:I
*+ wbs_stb_i:I wbs_cyc_i:I wbs_we_i:I wbs_sel_i[3:0]:I wbs_dat_i[31:0]:I wbs_adr_i[31:0]:I wbs_ack_o:O
*+ wbs_dat_o[31:0]:O la_data_in[127:0]:I la_data_out[127:0]:O io_in[26:0]:I io_in_3v3[26:0]:I user_clock2:I
*+ io_out[26:0]:O io_oeb[26:0]:O gpio_analog[17:0]:B gpio_noesd[17:0]:B io_analog[10:0]:B io_clamp_high[2:0]:B
*+ io_clamp_low[2:0]:B user_irq[2:0]:O la_oenb[127:0]:I
x1 io_analog[10] vccd1 vdda1 io_analog[1] io_analog[2] io_analog[3] io_analog[4] vssd1 io_analog[5]
+ vdda2 vccd2 vssd1 vccd1 io_analog[5] vdda2 wbs_we_i vssd1 vccd2 wbs_we_i vccd2 wbs_we_i vdda1
+ wishbone_address_bus[31] wishbone_address_bus[30] wishbone_address_bus[29] wishbone_address_bus[28] wishbone_address_bus[27]
+ wishbone_address_bus[26] wishbone_address_bus[25] wishbone_address_bus[24] wishbone_address_bus[23] wishbone_address_bus[22]
+ wishbone_address_bus[21] wishbone_address_bus[20] wishbone_address_bus[19] wishbone_address_bus[18] wishbone_address_bus[17]
+ wishbone_address_bus[16] wishbone_address_bus[15] wishbone_address_bus[14] wishbone_address_bus[13] wishbone_address_bus[12]
+ wishbone_address_bus[11] wishbone_address_bus[10] wishbone_address_bus[9] wishbone_address_bus[8] wishbone_address_bus[7]
+ wishbone_address_bus[6] wishbone_address_bus[5] wishbone_address_bus[4] wishbone_address_bus[3] wishbone_address_bus[2]
+ wishbone_address_bus[1] wishbone_address_bus[0] CSA[15] CSA[14] CSA[13] CSA[12] CSA[11] CSA[10] CSA[9] CSA[8] CSA[7] CSA[6]
+ CSA[5] CSA[4] CSA[3] CSA[2] CSA[1] CSA[0] io_analog[0] wbs_dat_i[31] wbs_dat_i[30] wbs_dat_i[29]
+ wbs_dat_i[28] wbs_dat_i[27] wbs_dat_i[26] wbs_dat_i[25] wbs_dat_i[24] wbs_dat_i[23] wbs_dat_i[22] wbs_dat_i[21]
+ wbs_dat_i[20] wbs_dat_i[19] wbs_dat_i[18] wbs_dat_i[17] wbs_dat_i[16] wbs_dat_i[15] wbs_dat_i[14] wbs_dat_i[13]
+ wbs_dat_i[12] wbs_dat_i[11] wbs_dat_i[10] wbs_dat_i[9] wbs_dat_i[8] wbs_dat_i[7] wbs_dat_i[6] wbs_dat_i[5]
+ wbs_dat_i[4] wbs_dat_i[3] wbs_dat_i[2] wbs_dat_i[1] wbs_dat_i[0] gpio_analog[2] __UNCONNECTED_PIN__0 vssd1
+ gpio_analog[1] vccd1 wb_rst_i gpio_analog[0] __UNCONNECTED_PIN__1 wbs_dat_o[31] wbs_dat_o[30] wbs_dat_o[29]
+ wbs_dat_o[28] wbs_dat_o[27] wbs_dat_o[26] wbs_dat_o[25] wbs_dat_o[24] wbs_dat_o[23] wbs_dat_o[22] wbs_dat_o[21]
+ wbs_dat_o[20] wbs_dat_o[19] wbs_dat_o[18] wbs_dat_o[17] wbs_dat_o[16] wbs_dat_o[15] wbs_dat_o[14] wbs_dat_o[13]
+ wbs_dat_o[12] wbs_dat_o[11] wbs_dat_o[10] wbs_dat_o[9] wbs_dat_o[8] wbs_dat_o[7] wbs_dat_o[6] wbs_dat_o[5]
+ wbs_dat_o[4] wbs_dat_o[3] wbs_dat_o[2] wbs_dat_o[1] wbs_dat_o[0] wb_clk_i top_wrapper
.ends

* expanding   symbol:  RRAM_IMC/xschem/top_wrapper.sym # of pins=36
** sym_path: /home/nvm_user4/RRAM_IMC/xschem/top_wrapper.sym
** sch_path: /home/nvm_user4/RRAM_IMC/xschem/top_wrapper.sch
.subckt top_wrapper  SL VDD_LOW VDD_HIGH REF_CSA V2_REF_ADC V1_REF_ADC V0_REF_ADC V4_BL V3_BL V2_BL
+ V1_BL V4_SL V3_SL V2_SL V1_SL rd_sync_fifo_output_buffer_CSA V4_WL V3_WL rd_sync_fifo_output_buffer_ADC
+ V2_WL wbs_we_i V1_WL wishbone_address_bus[31] wishbone_address_bus[30] wishbone_address_bus[29]
+ wishbone_address_bus[28] wishbone_address_bus[27] wishbone_address_bus[26] wishbone_address_bus[25] wishbone_address_bus[24]
+ wishbone_address_bus[23] wishbone_address_bus[22] wishbone_address_bus[21] wishbone_address_bus[20] wishbone_address_bus[19]
+ wishbone_address_bus[18] wishbone_address_bus[17] wishbone_address_bus[16] wishbone_address_bus[15] wishbone_address_bus[14]
+ wishbone_address_bus[13] wishbone_address_bus[12] wishbone_address_bus[11] wishbone_address_bus[10] wishbone_address_bus[9]
+ wishbone_address_bus[8] wishbone_address_bus[7] wishbone_address_bus[6] wishbone_address_bus[5] wishbone_address_bus[4]
+ wishbone_address_bus[3] wishbone_address_bus[2] wishbone_address_bus[1] wishbone_address_bus[0] CSA[15] CSA[14] CSA[13]
+ CSA[12] CSA[11] CSA[10] CSA[9] CSA[8] CSA[7] CSA[6] CSA[5] CSA[4] CSA[3] CSA[2] CSA[1] CSA[0] VDD_PRE
+ wishbone_data_in[31] wishbone_data_in[30] wishbone_data_in[29] wishbone_data_in[28] wishbone_data_in[27]
+ wishbone_data_in[26] wishbone_data_in[25] wishbone_data_in[24] wishbone_data_in[23] wishbone_data_in[22]
+ wishbone_data_in[21] wishbone_data_in[20] wishbone_data_in[19] wishbone_data_in[18] wishbone_data_in[17]
+ wishbone_data_in[16] wishbone_data_in[15] wishbone_data_in[14] wishbone_data_in[13] wishbone_data_in[12]
+ wishbone_data_in[11] wishbone_data_in[10] wishbone_data_in[9] wishbone_data_in[8] wishbone_data_in[7]
+ wishbone_data_in[6] wishbone_data_in[5] wishbone_data_in[4] wishbone_data_in[3] wishbone_data_in[2] wishbone_data_in[1]
+ wishbone_data_in[0] ADC_OUT2[8] start_operation VSS ADC_OUT1[8] vdd1v8 rst ADC_OUT0[8] vdd3v3 wishbone_data_out[31]
+ wishbone_data_out[30] wishbone_data_out[29] wishbone_data_out[28] wishbone_data_out[27] wishbone_data_out[26]
+ wishbone_data_out[25] wishbone_data_out[24] wishbone_data_out[23] wishbone_data_out[22] wishbone_data_out[21]
+ wishbone_data_out[20] wishbone_data_out[19] wishbone_data_out[18] wishbone_data_out[17] wishbone_data_out[16]
+ wishbone_data_out[15] wishbone_data_out[14] wishbone_data_out[13] wishbone_data_out[12] wishbone_data_out[11]
+ wishbone_data_out[10] wishbone_data_out[9] wishbone_data_out[8] wishbone_data_out[7] wishbone_data_out[6]
+ wishbone_data_out[5] wishbone_data_out[4] wishbone_data_out[3] wishbone_data_out[2] wishbone_data_out[1]
+ wishbone_data_out[0] clk
*.PININFO clk:I rst:I vdd3v3:B wishbone_data_out[31:0]:O ADC_OUT0[8]:O vdd1v8:B start_operation:I
*+ wishbone_data_in[31:0]:I wishbone_address_bus[31:0]:I wbs_we_i:I VSS:B VDD_PRE:B V1_WL:B V2_WL:B V3_WL:B V4_WL:B V1_SL:B
*+ V2_SL:B V3_SL:B V4_SL:B V1_BL:B V2_BL:B V3_BL:B V4_BL:B V0_REF_ADC:B V1_REF_ADC:B V2_REF_ADC:B REF_CSA:B
*+ ADC_OUT1[8]:O ADC_OUT2[8]:O CSA[15:0]:O rd_sync_fifo_output_buffer_ADC:I rd_sync_fifo_output_buffer_CSA:I
*+ VDD_HIGH:B VDD_LOW:B SL:B
x1 SAEN_CSA REF_CSA CLK_EN_ADC[1] CLK_EN_ADC[0] PRE V2_REF_ADC V1_REF_ADC V0_REF_ADC ENABLE_CSA
+ IN0_BL[15] IN0_BL[14] IN0_BL[13] IN0_BL[12] IN0_BL[11] IN0_BL[10] IN0_BL[9] IN0_BL[8] IN0_BL[7] IN0_BL[6]
+ IN0_BL[5] IN0_BL[4] IN0_BL[3] IN0_BL[2] IN0_BL[1] IN0_BL[0] IN1_BL[15] IN1_BL[14] IN1_BL[13] IN1_BL[12]
+ IN1_BL[11] IN1_BL[10] IN1_BL[9] IN1_BL[8] IN1_BL[7] IN1_BL[6] IN1_BL[5] IN1_BL[4] IN1_BL[3] IN1_BL[2]
+ IN1_BL[1] IN1_BL[0] V4_BL V3_BL V2_BL V1_BL ENABLE_BL IN0_SL[15] IN0_SL[14] IN0_SL[13] IN0_SL[12] IN0_SL[11]
+ IN0_SL[10] IN0_SL[9] IN0_SL[8] IN0_SL[7] IN0_SL[6] IN0_SL[5] IN0_SL[4] IN0_SL[3] IN0_SL[2] IN0_SL[1] IN0_SL[0]
+ IN1_SL[15] IN1_SL[14] IN1_SL[13] IN1_SL[12] IN1_SL[11] IN1_SL[10] IN1_SL[9] IN1_SL[8] IN1_SL[7] IN1_SL[6]
+ IN1_SL[5] IN1_SL[4] IN1_SL[3] IN1_SL[2] IN1_SL[1] IN1_SL[0] V4_SL V3_SL V2_SL V1_SL ENABLE_SL IN0_WL[15]
+ IN0_WL[14] IN0_WL[13] IN0_WL[12] IN0_WL[11] IN0_WL[10] IN0_WL[9] IN0_WL[8] IN0_WL[7] IN0_WL[6] IN0_WL[5]
+ IN0_WL[4] IN0_WL[3] IN0_WL[2] IN0_WL[1] IN0_WL[0] IN1_WL[15] IN1_WL[14] IN1_WL[13] IN1_WL[12] IN1_WL[11]
+ IN1_WL[10] IN1_WL[9] IN1_WL[8] IN1_WL[7] IN1_WL[6] IN1_WL[5] IN1_WL[4] IN1_WL[3] IN1_WL[2] IN1_WL[1] IN1_WL[0]
+ V4_WL SL V3_WL VDD_PRE ADC_OUT2[15] ADC_OUT2[14] ADC_OUT2[13] ADC_OUT2[12] ADC_OUT2[11] ADC_OUT2[10]
+ ADC_OUT2[9] ADC_OUT2[8] ADC_OUT2[7] ADC_OUT2[6] ADC_OUT2[5] ADC_OUT2[4] ADC_OUT2[3] ADC_OUT2[2] ADC_OUT2[1]
+ ADC_OUT2[0] V2_WL ADC_OUT1[15] ADC_OUT1[14] ADC_OUT1[13] ADC_OUT1[12] ADC_OUT1[11] ADC_OUT1[10] ADC_OUT1[9]
+ ADC_OUT1[8] ADC_OUT1[7] ADC_OUT1[6] ADC_OUT1[5] ADC_OUT1[4] ADC_OUT1[3] ADC_OUT1[2] ADC_OUT1[1] ADC_OUT1[0] VSS
+ V1_WL ADC_OUT0[15] ADC_OUT0[14] ADC_OUT0[13] ADC_OUT0[12] ADC_OUT0[11] ADC_OUT0[10] ADC_OUT0[9]
+ ADC_OUT0[8] ADC_OUT0[7] ADC_OUT0[6] ADC_OUT0[5] ADC_OUT0[4] ADC_OUT0[3] ADC_OUT0[2] ADC_OUT0[1] ADC_OUT0[0]
+ VDD_LOW CSA[15] CSA[14] CSA[13] CSA[12] CSA[11] CSA[10] CSA[9] CSA[8] CSA[7] CSA[6] CSA[5] CSA[4] CSA[3]
+ CSA[2] CSA[1] CSA[0] ENABLE_WL VDD_HIGH RRAM_ANALOG
x2 rd_sync_fifo_output_buffer_CSA rd_sync_fifo_output_buffer_ADC ENABLE_CSA IN1_SL[15] IN1_SL[14]
+ IN1_SL[13] IN1_SL[12] IN1_SL[11] IN1_SL[10] IN1_SL[9] IN1_SL[8] IN1_SL[7] IN1_SL[6] IN1_SL[5] IN1_SL[4]
+ IN1_SL[3] IN1_SL[2] IN1_SL[1] IN1_SL[0] IN0_SL[15] IN0_SL[14] IN0_SL[13] IN0_SL[12] IN0_SL[11] IN0_SL[10]
+ IN0_SL[9] IN0_SL[8] IN0_SL[7] IN0_SL[6] IN0_SL[5] IN0_SL[4] IN0_SL[3] IN0_SL[2] IN0_SL[1] IN0_SL[0]
+ ADC_OUT2[15] ADC_OUT2[14] ADC_OUT2[13] ADC_OUT2[12] ADC_OUT2[11] ADC_OUT2[10] ADC_OUT2[9] ADC_OUT2[8]
+ ADC_OUT2[7] ADC_OUT2[6] ADC_OUT2[5] ADC_OUT2[4] ADC_OUT2[3] ADC_OUT2[2] ADC_OUT2[1] ADC_OUT2[0] IN1_BL[15]
+ IN1_BL[14] IN1_BL[13] IN1_BL[12] IN1_BL[11] IN1_BL[10] IN1_BL[9] IN1_BL[8] IN1_BL[7] IN1_BL[6] IN1_BL[5]
+ IN1_BL[4] IN1_BL[3] IN1_BL[2] IN1_BL[1] IN1_BL[0] ADC_OUT1[15] ADC_OUT1[14] ADC_OUT1[13] ADC_OUT1[12]
+ ADC_OUT1[11] ADC_OUT1[10] ADC_OUT1[9] ADC_OUT1[8] ADC_OUT1[7] ADC_OUT1[6] ADC_OUT1[5] ADC_OUT1[4] ADC_OUT1[3]
+ ADC_OUT1[2] ADC_OUT1[1] ADC_OUT1[0] IN0_BL[15] IN0_BL[14] IN0_BL[13] IN0_BL[12] IN0_BL[11] IN0_BL[10] IN0_BL[9]
+ IN0_BL[8] IN0_BL[7] IN0_BL[6] IN0_BL[5] IN0_BL[4] IN0_BL[3] IN0_BL[2] IN0_BL[1] IN0_BL[0] ADC_OUT0[15]
+ ADC_OUT0[14] ADC_OUT0[13] ADC_OUT0[12] ADC_OUT0[11] ADC_OUT0[10] ADC_OUT0[9] ADC_OUT0[8] ADC_OUT0[7] ADC_OUT0[6]
+ ADC_OUT0[5] ADC_OUT0[4] ADC_OUT0[3] ADC_OUT0[2] ADC_OUT0[1] ADC_OUT0[0] IN1_WL[15] IN1_WL[14] IN1_WL[13]
+ IN1_WL[12] IN1_WL[11] IN1_WL[10] IN1_WL[9] IN1_WL[8] IN1_WL[7] IN1_WL[6] IN1_WL[5] IN1_WL[4] IN1_WL[3]
+ IN1_WL[2] IN1_WL[1] IN1_WL[0] IN0_WL[15] IN0_WL[14] IN0_WL[13] IN0_WL[12] IN0_WL[11] IN0_WL[10] IN0_WL[9]
+ IN0_WL[8] IN0_WL[7] IN0_WL[6] IN0_WL[5] IN0_WL[4] IN0_WL[3] IN0_WL[2] IN0_WL[1] IN0_WL[0] CSA[15] CSA[14]
+ CSA[13] CSA[12] CSA[11] CSA[10] CSA[9] CSA[8] CSA[7] CSA[6] CSA[5] CSA[4] CSA[3] CSA[2] CSA[1] CSA[0]
+ SAEN_CSA wbs_we_i CLK_EN_ADC[1] CLK_EN_ADC[0] wishbone_address_bus[31] wishbone_address_bus[30]
+ wishbone_address_bus[29] wishbone_address_bus[28] wishbone_address_bus[27] wishbone_address_bus[26] wishbone_address_bus[25]
+ wishbone_address_bus[24] wishbone_address_bus[23] wishbone_address_bus[22] wishbone_address_bus[21] wishbone_address_bus[20]
+ wishbone_address_bus[19] wishbone_address_bus[18] wishbone_address_bus[17] wishbone_address_bus[16] wishbone_address_bus[15]
+ wishbone_address_bus[14] wishbone_address_bus[13] wishbone_address_bus[12] wishbone_address_bus[11] wishbone_address_bus[10]
+ wishbone_address_bus[9] wishbone_address_bus[8] wishbone_address_bus[7] wishbone_address_bus[6] wishbone_address_bus[5]
+ wishbone_address_bus[4] wishbone_address_bus[3] wishbone_address_bus[2] wishbone_address_bus[1] wishbone_address_bus[0] PRE
+ wishbone_data_in[31] wishbone_data_in[30] wishbone_data_in[29] wishbone_data_in[28] wishbone_data_in[27]
+ wishbone_data_in[26] wishbone_data_in[25] wishbone_data_in[24] wishbone_data_in[23] wishbone_data_in[22]
+ wishbone_data_in[21] wishbone_data_in[20] wishbone_data_in[19] wishbone_data_in[18] wishbone_data_in[17]
+ wishbone_data_in[16] wishbone_data_in[15] wishbone_data_in[14] wishbone_data_in[13] wishbone_data_in[12]
+ wishbone_data_in[11] wishbone_data_in[10] wishbone_data_in[9] wishbone_data_in[8] wishbone_data_in[7]
+ wishbone_data_in[6] wishbone_data_in[5] wishbone_data_in[4] wishbone_data_in[3] wishbone_data_in[2] wishbone_data_in[1]
+ wishbone_data_in[0] COL_SELECT ENABLE_BL start_operation vdd3v3 ENABLE_SL vdd1v8 rst ENABLE_WL VSS
+ wishbone_data_out[31] wishbone_data_out[30] wishbone_data_out[29] wishbone_data_out[28] wishbone_data_out[27]
+ wishbone_data_out[26] wishbone_data_out[25] wishbone_data_out[24] wishbone_data_out[23] wishbone_data_out[22]
+ wishbone_data_out[21] wishbone_data_out[20] wishbone_data_out[19] wishbone_data_out[18] wishbone_data_out[17]
+ wishbone_data_out[16] wishbone_data_out[15] wishbone_data_out[14] wishbone_data_out[13] wishbone_data_out[12]
+ wishbone_data_out[11] wishbone_data_out[10] wishbone_data_out[9] wishbone_data_out[8] wishbone_data_out[7]
+ wishbone_data_out[6] wishbone_data_out[5] wishbone_data_out[4] wishbone_data_out[3] wishbone_data_out[2]
+ wishbone_data_out[1] wishbone_data_out[0] clk RRAM_CONTROLLER
.ends


* expanding   symbol:  RRAM_IMC/xschem/RRAM_ANALOG.sym # of pins=38
** sym_path: /home/nvm_user4/RRAM_IMC/xschem/RRAM_ANALOG.sym
** sch_path: /home/nvm_user4/RRAM_IMC/xschem/RRAM_ANALOG.sch
.subckt RRAM_ANALOG  SAEN_CSA REF_CSA CLK_EN_ADC[1] CLK_EN_ADC[0] PRE V2_REF_ADC V1_REF_ADC
+ V0_REF_ADC ENABLE_CSA IN0_BL[15] IN0_BL[14] IN0_BL[13] IN0_BL[12] IN0_BL[11] IN0_BL[10] IN0_BL[9] IN0_BL[8]
+ IN0_BL[7] IN0_BL[6] IN0_BL[5] IN0_BL[4] IN0_BL[3] IN0_BL[2] IN0_BL[1] IN0_BL[0] IN1_BL[15] IN1_BL[14]
+ IN1_BL[13] IN1_BL[12] IN1_BL[11] IN1_BL[10] IN1_BL[9] IN1_BL[8] IN1_BL[7] IN1_BL[6] IN1_BL[5] IN1_BL[4]
+ IN1_BL[3] IN1_BL[2] IN1_BL[1] IN1_BL[0] V4_BL V3_BL V2_BL V1_BL ENABLE_BL IN0_SL[15] IN0_SL[14] IN0_SL[13]
+ IN0_SL[12] IN0_SL[11] IN0_SL[10] IN0_SL[9] IN0_SL[8] IN0_SL[7] IN0_SL[6] IN0_SL[5] IN0_SL[4] IN0_SL[3]
+ IN0_SL[2] IN0_SL[1] IN0_SL[0] IN1_SL[15] IN1_SL[14] IN1_SL[13] IN1_SL[12] IN1_SL[11] IN1_SL[10] IN1_SL[9]
+ IN1_SL[8] IN1_SL[7] IN1_SL[6] IN1_SL[5] IN1_SL[4] IN1_SL[3] IN1_SL[2] IN1_SL[1] IN1_SL[0] V4_SL V3_SL V2_SL
+ V1_SL ENABLE_SL IN0_WL[15] IN0_WL[14] IN0_WL[13] IN0_WL[12] IN0_WL[11] IN0_WL[10] IN0_WL[9] IN0_WL[8]
+ IN0_WL[7] IN0_WL[6] IN0_WL[5] IN0_WL[4] IN0_WL[3] IN0_WL[2] IN0_WL[1] IN0_WL[0] IN1_WL[15] IN1_WL[14]
+ IN1_WL[13] IN1_WL[12] IN1_WL[11] IN1_WL[10] IN1_WL[9] IN1_WL[8] IN1_WL[7] IN1_WL[6] IN1_WL[5] IN1_WL[4]
+ IN1_WL[3] IN1_WL[2] IN1_WL[1] IN1_WL[0] V4_WL SL V3_WL VDD_PRE ADC_OUT2[15] ADC_OUT2[14] ADC_OUT2[13]
+ ADC_OUT2[12] ADC_OUT2[11] ADC_OUT2[10] ADC_OUT2[9] ADC_OUT2[8] ADC_OUT2[7] ADC_OUT2[6] ADC_OUT2[5] ADC_OUT2[4]
+ ADC_OUT2[3] ADC_OUT2[2] ADC_OUT2[1] ADC_OUT2[0] V2_WL ADC_OUT1[15] ADC_OUT1[14] ADC_OUT1[13] ADC_OUT1[12]
+ ADC_OUT1[11] ADC_OUT1[10] ADC_OUT1[9] ADC_OUT1[8] ADC_OUT1[7] ADC_OUT1[6] ADC_OUT1[5] ADC_OUT1[4] ADC_OUT1[3]
+ ADC_OUT1[2] ADC_OUT1[1] ADC_OUT1[0] VSS V1_WL ADC_OUT0[15] ADC_OUT0[14] ADC_OUT0[13] ADC_OUT0[12] ADC_OUT0[11]
+ ADC_OUT0[10] ADC_OUT0[9] ADC_OUT0[8] ADC_OUT0[7] ADC_OUT0[6] ADC_OUT0[5] ADC_OUT0[4] ADC_OUT0[3] ADC_OUT0[2]
+ ADC_OUT0[1] ADC_OUT0[0] VDD_LOW CSA[15] CSA[14] CSA[13] CSA[12] CSA[11] CSA[10] CSA[9] CSA[8] CSA[7] CSA[6]
+ CSA[5] CSA[4] CSA[3] CSA[2] CSA[1] CSA[0] ENABLE_WL VDD_HIGH
*.PININFO VDD_HIGH:B VDD_LOW:B CSA[15:0]:O V1_WL:I V2_WL:I V3_WL:I V4_WL:I IN1_WL[15:0]:I
*+ IN0_WL[15:0]:I ENABLE_SL:I V1_SL:I V2_SL:I V3_SL:I V4_SL:I IN1_SL[15:0]:I IN0_SL[15:0]:I ENABLE_BL:I V1_BL:I
*+ V2_BL:I V3_BL:I V4_BL:I IN1_BL[15:0]:I IN0_BL[15:0]:I ENABLE_CSA:I V0_REF_ADC:I V1_REF_ADC:I V2_REF_ADC:I
*+ PRE:I VSS:B ADC_OUT0[15:0]:O ADC_OUT1[15:0]:O ADC_OUT2[15:0]:O CLK_EN_ADC[1:0]:I REF_CSA:I SAEN_CSA:I
*+ ENABLE_WL:I VDD_PRE:B SL:B
.ends


* expanding   symbol:  RRAM_IMC/xschem/RRAM_CONTROLLER.sym # of pins=30
** sym_path: /home/nvm_user4/RRAM_IMC/xschem/RRAM_CONTROLLER.sym
** sch_path: /home/nvm_user4/RRAM_IMC/xschem/RRAM_CONTROLLER.sch
.subckt RRAM_CONTROLLER  rd_sync_fifo_output_buffer_CSA rd_sync_fifo_output_buffer_ADC ENABLE_CSA
+ IN1_SL[15] IN1_SL[14] IN1_SL[13] IN1_SL[12] IN1_SL[11] IN1_SL[10] IN1_SL[9] IN1_SL[8] IN1_SL[7] IN1_SL[6]
+ IN1_SL[5] IN1_SL[4] IN1_SL[3] IN1_SL[2] IN1_SL[1] IN1_SL[0] IN0_SL[15] IN0_SL[14] IN0_SL[13] IN0_SL[12]
+ IN0_SL[11] IN0_SL[10] IN0_SL[9] IN0_SL[8] IN0_SL[7] IN0_SL[6] IN0_SL[5] IN0_SL[4] IN0_SL[3] IN0_SL[2]
+ IN0_SL[1] IN0_SL[0] ADC_OUT2[15] ADC_OUT2[14] ADC_OUT2[13] ADC_OUT2[12] ADC_OUT2[11] ADC_OUT2[10] ADC_OUT2[9]
+ ADC_OUT2[8] ADC_OUT2[7] ADC_OUT2[6] ADC_OUT2[5] ADC_OUT2[4] ADC_OUT2[3] ADC_OUT2[2] ADC_OUT2[1] ADC_OUT2[0]
+ IN1_BL[15] IN1_BL[14] IN1_BL[13] IN1_BL[12] IN1_BL[11] IN1_BL[10] IN1_BL[9] IN1_BL[8] IN1_BL[7] IN1_BL[6]
+ IN1_BL[5] IN1_BL[4] IN1_BL[3] IN1_BL[2] IN1_BL[1] IN1_BL[0] ADC_OUT1[15] ADC_OUT1[14] ADC_OUT1[13]
+ ADC_OUT1[12] ADC_OUT1[11] ADC_OUT1[10] ADC_OUT1[9] ADC_OUT1[8] ADC_OUT1[7] ADC_OUT1[6] ADC_OUT1[5] ADC_OUT1[4]
+ ADC_OUT1[3] ADC_OUT1[2] ADC_OUT1[1] ADC_OUT1[0] IN0_BL[15] IN0_BL[14] IN0_BL[13] IN0_BL[12] IN0_BL[11]
+ IN0_BL[10] IN0_BL[9] IN0_BL[8] IN0_BL[7] IN0_BL[6] IN0_BL[5] IN0_BL[4] IN0_BL[3] IN0_BL[2] IN0_BL[1] IN0_BL[0]
+ ADC_OUT0[15] ADC_OUT0[14] ADC_OUT0[13] ADC_OUT0[12] ADC_OUT0[11] ADC_OUT0[10] ADC_OUT0[9] ADC_OUT0[8]
+ ADC_OUT0[7] ADC_OUT0[6] ADC_OUT0[5] ADC_OUT0[4] ADC_OUT0[3] ADC_OUT0[2] ADC_OUT0[1] ADC_OUT0[0] IN1_WL[15]
+ IN1_WL[14] IN1_WL[13] IN1_WL[12] IN1_WL[11] IN1_WL[10] IN1_WL[9] IN1_WL[8] IN1_WL[7] IN1_WL[6] IN1_WL[5]
+ IN1_WL[4] IN1_WL[3] IN1_WL[2] IN1_WL[1] IN1_WL[0] IN0_WL[15] IN0_WL[14] IN0_WL[13] IN0_WL[12] IN0_WL[11]
+ IN0_WL[10] IN0_WL[9] IN0_WL[8] IN0_WL[7] IN0_WL[6] IN0_WL[5] IN0_WL[4] IN0_WL[3] IN0_WL[2] IN0_WL[1] IN0_WL[0]
+ CSA[15] CSA[14] CSA[13] CSA[12] CSA[11] CSA[10] CSA[9] CSA[8] CSA[7] CSA[6] CSA[5] CSA[4] CSA[3] CSA[2]
+ CSA[1] CSA[0] SAEN_CSA wbs_we_i CLK_EN_ADC[1] CLK_EN_ADC[0] wishbone_address_bus[31]
+ wishbone_address_bus[30] wishbone_address_bus[29] wishbone_address_bus[28] wishbone_address_bus[27] wishbone_address_bus[26]
+ wishbone_address_bus[25] wishbone_address_bus[24] wishbone_address_bus[23] wishbone_address_bus[22] wishbone_address_bus[21]
+ wishbone_address_bus[20] wishbone_address_bus[19] wishbone_address_bus[18] wishbone_address_bus[17] wishbone_address_bus[16]
+ wishbone_address_bus[15] wishbone_address_bus[14] wishbone_address_bus[13] wishbone_address_bus[12] wishbone_address_bus[11]
+ wishbone_address_bus[10] wishbone_address_bus[9] wishbone_address_bus[8] wishbone_address_bus[7] wishbone_address_bus[6]
+ wishbone_address_bus[5] wishbone_address_bus[4] wishbone_address_bus[3] wishbone_address_bus[2] wishbone_address_bus[1]
+ wishbone_address_bus[0] PRE wishbone_data_in[31] wishbone_data_in[30] wishbone_data_in[29] wishbone_data_in[28]
+ wishbone_data_in[27] wishbone_data_in[26] wishbone_data_in[25] wishbone_data_in[24] wishbone_data_in[23]
+ wishbone_data_in[22] wishbone_data_in[21] wishbone_data_in[20] wishbone_data_in[19] wishbone_data_in[18]
+ wishbone_data_in[17] wishbone_data_in[16] wishbone_data_in[15] wishbone_data_in[14] wishbone_data_in[13]
+ wishbone_data_in[12] wishbone_data_in[11] wishbone_data_in[10] wishbone_data_in[9] wishbone_data_in[8]
+ wishbone_data_in[7] wishbone_data_in[6] wishbone_data_in[5] wishbone_data_in[4] wishbone_data_in[3] wishbone_data_in[2]
+ wishbone_data_in[1] wishbone_data_in[0] COL_SELECT ENABLE_BL start_operation vdd3v3 ENABLE_SL vdd1v8 rst ENABLE_WL VSS
+ wishbone_data_out[31] wishbone_data_out[30] wishbone_data_out[29] wishbone_data_out[28] wishbone_data_out[27]
+ wishbone_data_out[26] wishbone_data_out[25] wishbone_data_out[24] wishbone_data_out[23] wishbone_data_out[22]
+ wishbone_data_out[21] wishbone_data_out[20] wishbone_data_out[19] wishbone_data_out[18] wishbone_data_out[17]
+ wishbone_data_out[16] wishbone_data_out[15] wishbone_data_out[14] wishbone_data_out[13] wishbone_data_out[12]
+ wishbone_data_out[11] wishbone_data_out[10] wishbone_data_out[9] wishbone_data_out[8] wishbone_data_out[7]
+ wishbone_data_out[6] wishbone_data_out[5] wishbone_data_out[4] wishbone_data_out[3] wishbone_data_out[2]
+ wishbone_data_out[1] wishbone_data_out[0] clk
*.PININFO clk:I rst:I VSS:B wishbone_data_out[31:0]:O ENABLE_WL:O start_operation:I
*+ wishbone_data_in[31:0]:I wishbone_address_bus[31:0]:I wbs_we_i:I CSA[15:0]:I ADC_OUT0[15:0]:I ADC_OUT1[15:0]:I
*+ ADC_OUT2[15:0]:I ENABLE_CSA:I rd_sync_fifo_output_buffer_ADC:I rd_sync_fifo_output_buffer_CSA:I vdd1v8:B vdd3v3:B
*+ ENABLE_SL:O ENABLE_BL:O COL_SELECT:O PRE:O CLK_EN_ADC[1:0]:O SAEN_CSA:O IN0_WL[15:0]:O IN1_WL[15:0]:O
*+ IN0_BL[15:0]:O IN1_BL[15:0]:O IN0_SL[15:0]:O IN1_SL[15:0]:O
.ends

.end
